module vecs

pub struct Physics {
	pub mut:
	x_speed f64
	y_speed f64
}