module vecs

pub struct Gravity {
}
