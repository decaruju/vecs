module vecs

interface Component {}
