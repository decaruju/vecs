module vecs

pub struct Position {
pub mut:
	x f64
	y f64
}
